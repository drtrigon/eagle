Ultra_RBBB_V01
C2 0 8 100nF IC=0
R1 1 5 220
C1 0 7 100nF IC=0
C3 4 5 100nF IC=0

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
